module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
		case (Address[9:2])
			8'd0:    Instruction <= 32'b00001000000000000000000000001110;
			8'd1:    Instruction <= 32'b00001000000000000000000000010011;
			8'd2:    Instruction <= 32'b00001000000000000000000000010011;
			8'd3:    Instruction <= 32'b00010000100001010000000000000011;
			8'd4:    Instruction <= 32'b00000000100001010100000000101010;
			8'd5:    Instruction <= 32'b00010001000100000000000000000011;
			8'd6:    Instruction <= 32'b00001000000000000000000000001011;
			8'd7:    Instruction <= 32'b00000000100000000001000000100000;
			8'd8:    Instruction <= 32'b00001000000000000000000000010011;
			8'd9:    Instruction <= 32'b00000000101001000010100000100010;
			8'd10:    Instruction <= 32'b00001000000000000000000000000011;
			8'd11:    Instruction <= 32'b00000000100001010010000000100010;
			8'd12:    Instruction <= 32'b00000000000000000000000000000000;
			8'd13:    Instruction <= 32'b00001000000000000000000000000011;
			8'd14:    Instruction <= 32'b00100000000001000000000001111101;
			8'd15:    Instruction <= 32'b00000000000000000000000000000000;
			8'd16:    Instruction <= 32'b00100000000001010000000000101000;
			8'd17:    Instruction <= 32'b00100000000100000000000000000001;
			8'd18:    Instruction <= 32'b00001000000000000000000000000011;
			8'd19:    Instruction <= 32'b00000000010000000001000000100000;			
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule