module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
		case (Address[9:2])
			8'd0: Instruction <= 32'b00001000000000000000000000001110;
8'd1: Instruction <= 32'b00001000000000000000000000100111;
8'd2: Instruction <= 32'b00001000000000000000000000100111;
8'd3: Instruction <= 32'b00010000100001010000000000000011;
8'd4: Instruction <= 32'b00000000100001010100000000101010;
8'd5: Instruction <= 32'b00010001000100000000000000000011;
8'd6: Instruction <= 32'b00001000000000000000000000001011;
8'd7: Instruction <= 32'b00000000100000000001000000100000;
8'd8: Instruction <= 32'b00001000000000000000000000100111;
8'd9: Instruction <= 32'b00000000101001000010100000100010;
8'd10: Instruction <= 32'b00001000000000000000000000000011;
8'd11: Instruction <= 32'b00000000100001010010000000100010;
8'd12: Instruction <= 32'b00000000000000000000000000000000;
8'd13: Instruction <= 32'b00001000000000000000000000000011;
8'd14: Instruction <= 32'b00111100000000010100000000000000;
8'd15: Instruction <= 32'b00110100001000010000000000100000;
8'd16: Instruction <= 32'b00000000000000010100000000100000;
8'd17: Instruction <= 32'b10001101000010010000000000000000;
8'd18: Instruction <= 32'b00110001001010010000000000001000;
8'd19: Instruction <= 32'b00010001001000001111111111111101;
8'd20: Instruction <= 32'b00000000000000000000000000000000;
8'd21: Instruction <= 32'b00111100000000010100000000000000;
8'd22: Instruction <= 32'b00110100001000010000000000011100;
8'd23: Instruction <= 32'b00000000000000010010000000100000;
8'd24: Instruction <= 32'b10001100100001000000000000000000;
8'd25: Instruction <= 32'b00000000000000000000000000000000;
8'd26: Instruction <= 32'b00111100000000010100000000000000;
8'd27: Instruction <= 32'b00110100001000010000000000100000;
8'd28: Instruction <= 32'b00000000000000010100000000100000;
8'd29: Instruction <= 32'b10001101000010010000000000000000;
8'd30: Instruction <= 32'b00110001001010010000000000001000;
8'd31: Instruction <= 32'b00010001001000001111111111111101;
8'd32: Instruction <= 32'b00000000000000000000000000000000;
8'd33: Instruction <= 32'b00111100000000010100000000000000;
8'd34: Instruction <= 32'b00110100001000010000000000011100;
8'd35: Instruction <= 32'b00000000000000010010100000100000;
8'd36: Instruction <= 32'b10001100101001010000000000000000;
8'd37: Instruction <= 32'b00100000000100000000000000000001;
8'd38: Instruction <= 32'b00001000000000000000000000000011;
8'd39: Instruction <= 32'b00000000010000000001000000100000;
8'd40: Instruction <= 32'b00111100000000010100000000000000;
8'd41: Instruction <= 32'b00110100001000010000000000011000;
8'd42: Instruction <= 32'b00000000000000010011000000100000;
8'd43: Instruction <= 32'b10101100110000100000000000000000;	
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule