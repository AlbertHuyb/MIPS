module Forward();


endmodule

module 