module IFIDReg();

endmodule // IFIDReg

module IDEXReg();

endmodule // IDEXReg

module EXMEMReg();

endmodule // EXMEMReg

module MEMWBReg();

endmodule // MEMWBReg