module BCD(
    din,
    dout
);
input   [3:0]   din;
output  [6:0]   dout;

assign  dout=(din==4'h0)?7'b1000000: //64
             (din==4'h1)?7'b1111001: //121
             (din==4'h2)?7'b0100100: //36
             (din==4'h3)?7'b0110000: //48
             (din==4'h4)?7'b0011001: //25
             (din==4'h5)?7'b0010010: //18
             (din==4'h6)?7'b0000010: //2
             (din==4'h7)?7'b1111000: //120
             (din==4'h8)?7'b0000000: //0
             (din==4'h9)?7'b0010000: //16
             (din==4'hA)?7'b0001000: //8
             (din==4'hB)?7'b0000011: //3
             (din==4'hC)?7'b1000110: //134
             (din==4'hD)?7'b0100001: //33
             (din==4'hE)?7'b0000110: //6
             (din==4'hF)?7'b0001110:7'b0; //14
endmodule