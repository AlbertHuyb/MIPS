/*
Write your code for reg between module here.
And add what you need.
Good Luck!
*/

module IFIDReg();

endmodule // IFIDReg

module IDEXReg();

endmodule // IDEXReg

module EXMEMReg();

endmodule // EXMEMReg

module MEMWBReg();

endmodule // MEMWBReg